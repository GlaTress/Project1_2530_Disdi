LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY twoComp IS
  GENERIC ( N : INTEGER := 4 );
  PORT (
    X : IN  STD_LOGIC_VECTOR(N-1 DOWNTO 0);
    Y : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE twoCompArch OF twoComp IS
  SIGNAL Aux : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
BEGIN

  Aux(0) <= '0';

  GEN_SEEN : FOR i IN 0 TO N-2 GENERATE
    Aux(i+1) <= Aux(i) OR X(i);
  END GENERATE;

  GEN_Y : FOR i IN 0 TO N-1 GENERATE
    Y(i)     <= X(i) XOR Aux(i);
  END GENERATE;

END ARCHITECTURE;
